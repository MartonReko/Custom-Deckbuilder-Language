//OUTDATED
Game{
    Name: xyz;
    Stages: [a,b,c];
    Player: c1;
}

Stage a{
    Length: 1;
    Max-width: 1;
    Min-width: 1;
    FillWith: [node1];
    MustContain: [3x node2];
    EndsWith: node3;
}

Node node1{
    Enemies: [
    2x enemy1,
    1x enemy2 or
    2x enemy1
    ];
    Rewards: [
		3x common with chance 50% or
		2x rare with chance 40% or
		6x common with chance 10%
    ];
}

Character c1{
    Health: 1;
    EffectEveryTurn: [];
}

Effect e1{
    Outgoing damage is damage * 2.2;
    Incoming damage is damage * 0.9;

    Deal 122 damage instantly to target
    Apply [e2,e3] for 6 turns to enemies
}

Card c1{
    Rarity: rarity1;
    ValidTargets: [self, enemies];
    Apply [e4,e5]
}