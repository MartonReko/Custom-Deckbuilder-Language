Game{
    Name: My_Wonderful_Game;
    Stages: [
    beginnerStage,
    advancedStage
    ];
    Player: MyCharacter;
}

Character MyCharacter{
    Health: 75;
    EffectEveryTurn: [smallHeal];
    Deck: [10x strike];
}

Effect smallHeal{
    Deal -1 damage instantly;
}

Stage beginnerStage{
    Length: 10;
    Length: 10;
    Max-width: 5;
    Min-width: 2;
    FillWith: [easyNode];
    MustContain: [1x eliteNode, 2x normalNode];
    EndsWith: bossNode;
}

Node eliteNode{
    Enemies: [1x  eliteEnemy];
    Rewards: [3x rare with chance 100%];
}

Stage advancedStage{
    Length: 5;
    Max-width: 3;
    Min-width: 1;
    FillWith: [easyNode,eliteNode];
    MustContain: [3x eliteNode];
    EndsWith: bossNode;
}

Node easyNode{
    Enemies: [
    2x easyEnemy
    ];
    Rewards: [
		3x common with chance 80%,
		2x rare with chance 20%
    ];
}
Node normalNode{
    Enemies: [
    3x easyEnemy
    ];
    Rewards: [
		3x common with chance 50%,
		2x rare with chance 50%
    ];
}



Node bossNode{
    Enemies: [
    1x bossEnemy
    ];
    Rewards: [
        3x rare with chance 100%
    ];
}

Enemy easyEnemy{
    Health: 10;
    Actions: [basicEnemyAttack player];
}

Enemy enemy_hard{
    Health: 30;
    Actions: [basicEnemyAttack player];
}

Enemy eliteEnemy{
    Health: 50;
    Actions: [basicEnemyAttack player,statusAttack player];
}


Enemy bossEnemy{
    Health: 100;
    Actions: [bossAttack player, 2x statusAttack player, bossBuff self];
}
EnemyAction bossAttack{
    Apply: [bossDamageEffect, poisonEffect];
}
EnemyAction statusAttack{
    Apply: [curseEffect, poisonEffect];
}
EnemyAction bossBuff{
    Apply: [bossBuffEffect];
}
Effect bossDamageEffect{
    Deal 20 damage instantly;
}
Effect bossBuffEffect{
    Outgoing damage is 1.25x;
    Incoming damage is 0.75x;
}

EnemyAction basicEnemyAttack{
    Apply: [2x basicAttack, poisonEffect];
}




Effect curseEffect{
    Outgoing damage is 0.75x;
    Incoming damage is 1.2x;
}
Card superCard{
    Rarity: rare;
    ValidTargets: [enemy];
    Apply: [10x basicAttack, 5x weakness, 2x poisonEffect];
}
Effect poisonEffect{
    Deal 3 damage end of turn;
}
Effect basicAttack{
    Deal baseDamage * 2 damage instantly;
}
Effect weakness{
    Outgoing damage is 0.75x;
}

int baseDamage = 5;

Card strike{
    Rarity: common;
    ValidTargets: [enemy];
    Apply: [basicAttack];
}
Card heal{
    Rarity: rare;
    ValidTargets: [player];
    Apply: [smallHeal];
}

Card poison{
    Rarity: common;
    ValidTargets: [player, enemy];
    Apply: [2x poisonEffect, weakness];
}