Game{
    Name: My_Wonderful_Game;
    Stages: [
    stage_beginner,
    stage_advanced
    ];
    Player: Bob;
}

Character Bob{
    Health: 75;
    EffectEveryTurn: [small_heal];
    Deck: [10x strike];
}

Effect small_heal{
    Deal -1 damage instantly;
}

Stage stage_beginner{
    Length: 3;
    Max-width: 3;
    Min-width: 1;
    FillWith: [node_easy];
    MustContain: [1x node_elite];
    EndsWith: node_boss;
}

Stage stage_advanced{
    Length: 5;
    Max-width: 3;
    Min-width: 1;
    FillWith: [node_easy,node_elite];
    MustContain: [3x node_elite];
    EndsWith: node_boss;
}

Node node_easy{
    Enemies: [
    2x enemy_easy
    ];
    Rewards: [
		3x rarity_common with chance 80%,
		2x rarity_rare with chance 20%
    ];
}

Node node_elite{
    Enemies: [
    1x  enemy_elite
    ];
    Rewards: [
        3x rarity_rare with chance 100%
    ];
}

Node node_boss{
    Enemies: [
    1x enemy_boss
    ];
    Rewards: [
        3x rarity_rare with chance 100%
    ];
}

Enemy enemy_easy{
    Health: 10;
    Actions: [basicAttack player];
}

Enemy enemy_hard{
    Health: 30;
    Actions: [basicAttack player];
}

Enemy enemy_elite{
    Health: 50;
    Actions: [basicAttack player,statusAttack player];
}

Enemy enemy_boss{
    Health: 100;
    Actions: [basicAttack player,3x statusAttack player];
}

EnemyAction basicAttack{
    Apply: [2x attack_basic, effect_poison];
}

EnemyAction statusAttack{
    Apply: [curse, effect_poison];
}

Effect attack_basic{
    Deal 5 damage instantly;
}

Effect curse{
    Outgoing damage is 0.75x;
    Incoming damage is 1.2x;
}

Effect effect_poison{
    Deal 3 damage end of turn;
}

Card strike{
    Rarity: rarity_common;
    ValidTargets: [enemy];
    Apply: [attack_basic];
}

Card heal{
    Rarity: rarity_rare;
    ValidTargets: [player];
    Apply: [small_heal];
}

Card poison{
    Rarity: rarity_common;
    ValidTargets: [player];
    Apply: [2x effect_poison];
}