Game{
    Name: My_Wonderful_Game;
    Stages: [
    stage_beginner,
    stage_advanced
    ];
    Player: ThePlayer;
}

Character The_Player{
    Health: 100;
    EffectEveryTurn: [miniscule_healing];
}

Stage stage_beginner{
    Length: 5;
    Max-width: 3;
    Min-width: 1;
    FillWith: [node_easy];
    MustContain: [1x node_elite];
    EndsWith: node_boss;
}

Stage stage_advanced{
    Length: 5;
    Max-width: 3;
    Min-width: 1;
    FillWith: [node_easy,node_elite];
    MustContain: [3x node_elite];
    EndsWith: node_boss;
}

Node node_easy{
    Enemies: [
    2x enemy_easy,
    1x enemy_hard or
    4x enemy_easy
    ];
    Rewards: [
		3x rarity_common with chance 80% or
		2x rarity_rare with chance 20%
    ];
}

Node node_elite{
    Enemies: [
    1x  enemy_elite
    ];
    Rewards: [
        3x rarity_rare with chance 100%
    ];
}

Node node_boss{
    Enemies: [
    1x enemy_boss or
    2x enemy_elite
    ];
    Rewards: [
        6x rarity_rare with chance 100%
    ];
}

Enemy enemy_easy{
    Health: 10;
    Actions: [attack_basic player];
}

Enemy enemy_hard{
    Health: 30;
    Actions: [attack_basic player];
}

Enemy enemy_elite{
    Health: 50;
    Actions: [attack_elite player, curse player];
}

Enemy enemy_boss{
    Health: 100;
    Actions: [attack_boss player, 2x curse player];
}

Effect attack_basic{
    Deal 5 damage instantly;
}

Effect attack_elite{
    Deal 15 damage instantly;
}

Effect curse{
    Outgoing damage is damage * 0.9;
    Incoming damage is damage * 1.2;
}

Effect strike_effect(int amount){
    Deal amount damage instantly;
}

// TODO
Effect effect_heal(int amount){
    Deal (-1 * amount) damage instantly;
}

Effect effect_poison(int amount){
    Deal amount damage end of turn;
}

Card strike{
    Rarity: rarity_common;
    ValidTargets: [enemy];
    Apply: [strike_effect(7)];
}

Card heal{
    Rarity: rarity_rare;
    ValidTargets: [player];
    Apply: [effect_heal(12)];
}

Card poison{
    Rarity: rarity_common;
    ValidTargets: [player];
    Apply: [2x effect_poison(2)];
}

int testInt = 5;
string testString = "asd";
double testDouble = 1.2;
bool testBoolean = false;